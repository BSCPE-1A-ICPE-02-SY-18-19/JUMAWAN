CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 52 187 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.89884e-315 0
0
2 +V
167 676 273 0 1 3
0 16
0
0 0 54256 180
3 10V
6 -2 27 6
3 V10
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9968 0 0
2
5.89884e-315 0
0
2 +V
167 531 269 0 1 3
0 17
0
0 0 54256 180
3 10V
6 -2 27 6
2 V9
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9281 0 0
2
5.89884e-315 0
0
2 +V
167 388 265 0 1 3
0 18
0
0 0 54256 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
5.89884e-315 0
0
2 +V
167 219 263 0 1 3
0 10
0
0 0 54256 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7168 0 0
2
5.89884e-315 0
0
2 +V
167 676 132 0 1 3
0 21
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3171 0 0
2
5.89884e-315 0
0
2 +V
167 531 133 0 1 3
0 22
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89884e-315 0
0
2 +V
167 386 126 0 1 3
0 23
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.89884e-315 0
0
7 Pulser~
4 89 303 0 10 12
0 25 26 19 27 0 0 5 5 5
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5283 0 0
2
5.89884e-315 0
0
9 2-In AND~
219 590 65 0 3 22
0 15 2 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6874 0 0
2
5.89884e-315 0
0
9 2-In AND~
219 397 56 0 3 22
0 12 13 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5305 0 0
2
5.89884e-315 0
0
9 CC 7-Seg~
183 912 78 0 18 19
10 9 8 7 6 5 4 3 28 29
0 0 0 1 1 0 1 2 2
0
0 0 21104 0
8 YELLOWCC
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
34 0 0
2
5.89884e-315 0
0
6 74LS48
188 849 200 0 14 29
0 11 2 13 12 30 31 3 4 5
6 7 8 9 32
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
969 0 0
2
5.89884e-315 0
0
6 74112~
219 676 224 0 7 32
0 21 14 19 14 16 33 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8402 0 0
2
5.89884e-315 0
0
6 74112~
219 531 224 0 7 32
0 22 15 19 15 17 34 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3751 0 0
2
5.89884e-315 0
0
6 74112~
219 386 224 0 7 32
0 23 12 19 12 18 35 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4292 0 0
2
5.89884e-315 0
0
6 74112~
219 219 223 0 7 32
0 24 20 19 20 10 36 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6118 0 0
2
5.89884e-315 0
0
2 +V
167 219 108 0 1 3
0 24
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
34 0 0
2
5.89884e-315 0
0
36
0 4 0 0 0 0 0 0 14 18 0 3
611 187
611 206
652 206
0 4 0 0 0 0 0 0 15 21 0 3
462 187
462 206
507 206
0 1 0 0 0 0 0 0 11 17 0 3
249 106
249 47
373 47
0 4 0 0 0 16 0 0 17 32 0 3
159 187
159 205
195 205
2 0 2 0 0 12416 0 13 0 0 19 4
817 173
761 173
761 88
562 88
7 7 3 0 0 4224 0 13 12 0 0 3
881 164
927 164
927 114
8 6 4 0 0 4224 0 13 12 0 0 3
881 173
921 173
921 114
9 5 5 0 0 4224 0 13 12 0 0 3
881 182
915 182
915 114
10 4 6 0 0 4224 0 13 12 0 0 3
881 191
909 191
909 114
11 3 7 0 0 4224 0 13 12 0 0 3
881 200
903 200
903 114
12 2 8 0 0 4224 0 13 12 0 0 3
881 209
897 209
897 114
13 1 9 0 0 4224 0 13 12 0 0 3
881 218
891 218
891 114
5 1 10 0 0 4224 0 17 5 0 0 2
219 235
219 248
7 1 11 0 0 12416 0 14 13 0 0 4
700 188
729 188
729 164
817 164
0 0 12 0 0 4096 0 0 0 17 0 2
739 106
743 106
0 3 13 0 0 4224 0 0 13 25 0 4
410 121
750 121
750 182
817 182
0 4 12 0 0 8320 0 0 13 27 0 5
249 188
249 106
739 106
739 191
817 191
3 2 14 0 0 4224 0 10 14 0 0 3
611 65
611 188
652 188
7 2 2 0 0 0 0 15 10 0 0 4
555 188
562 188
562 74
566 74
0 1 15 0 0 4096 0 0 10 21 0 2
462 56
566 56
3 2 15 0 0 0 0 11 15 0 0 4
418 56
462 56
462 188
507 188
5 1 16 0 0 4224 0 14 2 0 0 2
676 236
676 258
5 1 17 0 0 4224 0 15 3 0 0 2
531 236
531 254
5 1 18 0 0 8320 0 16 4 0 0 3
386 236
388 236
388 250
2 7 13 0 0 0 0 11 16 0 0 5
373 65
362 65
362 121
410 121
410 188
0 4 12 0 0 0 0 0 16 27 0 3
318 188
318 206
362 206
7 2 12 0 0 0 0 17 16 0 0 3
243 187
243 188
362 188
3 0 19 0 0 4096 0 17 0 0 31 2
189 196
189 294
3 0 19 0 0 0 0 16 0 0 31 2
356 197
356 294
3 0 19 0 0 0 0 15 0 0 31 2
501 197
501 294
3 3 19 0 0 4224 0 9 14 0 0 3
113 294
646 294
646 197
1 2 20 0 0 0 0 1 17 0 0 2
64 187
195 187
1 1 21 0 0 4224 0 6 14 0 0 2
676 141
676 161
1 1 22 0 0 4224 0 7 15 0 0 2
531 142
531 161
1 1 23 0 0 4224 0 8 16 0 0 2
386 135
386 161
1 1 24 0 0 4224 0 18 17 0 0 2
219 117
219 160
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
76 398 201 422
86 406 190 422
13 James Jumawan
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
